// fifo.v

// Generated using ACDS version 22.4 94

`timescale 1 ps / 1 ps
module fifo (
		input  wire [31:0] data,    //  fifo_input.datain
		input  wire        wrreq,   //            .wrreq
		input  wire        rdreq,   //            .rdreq
		input  wire        wrclk,   //            .wrclk
		input  wire        rdclk,   //            .rdclk
		input  wire        aclr,    //            .aclr
		output wire [31:0] q,       // fifo_output.dataout
		output wire        rdempty, //            .rdempty
		output wire        wrfull   //            .wrfull
	);

	fifo_fifo_1920_cgqugzq fifo_0 (
		.data    (data),    //   input,  width = 32,  fifo_input.datain
		.wrreq   (wrreq),   //   input,   width = 1,            .wrreq
		.rdreq   (rdreq),   //   input,   width = 1,            .rdreq
		.wrclk   (wrclk),   //   input,   width = 1,            .wrclk
		.rdclk   (rdclk),   //   input,   width = 1,            .rdclk
		.aclr    (aclr),    //   input,   width = 1,            .aclr
		.q       (q),       //  output,  width = 32, fifo_output.dataout
		.rdempty (rdempty), //  output,   width = 1,            .rdempty
		.wrfull  (wrfull)   //  output,   width = 1,            .wrfull
	);

endmodule
