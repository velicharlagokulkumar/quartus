module rom (
		output wire [31:0] q,       //       q.dataout
		input  wire [9:0]  address, // address.address
		input  wire        clock    //   clock.clk
	);
endmodule

