module golden_top (   
  input          FPGA_SYSTEM_CLK,
  input          FPGA_SYS_RESETN,
  input [7:0]    FPGA_SW,
  input [7:0]    FPGA_PB,
  output [7:0]   FPGA_LED_G,
  inout [15:0]   FPGA_GPIO,
  inout [12:0]   FPGA_TESTIO,
  inout          FPGA_TEST_ALERTN,
  
  input          REFCLK_GXPP0,
  input          REFCLK_GXPP2,
  input          REFCLK_GXEP0,
  input          REFCLK_GXEP1,
  input          REFCLK_GXEP2,
  input          REFCLK_GXEP3,   
  input          FPGA_GPIO_OUTCLKP,   
  input          FPGA_GPIO_REFCLKP0,   
  input          FPGA_GPIO_REFCLKP1,   
  input          FPGA_GPIO_REFCLKP2,   
  
  //I2C  
  inout          SODIMM_I2C_SDA,
  inout          SODIMM_I2C_SCL,
  inout          F2M_I2C_SCL,
  inout          F2M_I2C_SDA,
  inout          M2F_I2C_SCL,
  inout          M2F_I2C_SDA,
  inout          FPGA_TEST_SCL,
  inout          FPGA_TEST_SDA,
 
  //MXP		
  input  [3:0]   MXP_RXP,         
  input  [3:0]   MXP_RXN,         
  output [3:0]   MXP_TXP,         
  output [3:0]   MXP_TXN, 

  //ZQSFP		
  input  [3:0]   ZQSFP_RXP,         
  input  [3:0]   ZQSFP_RXN,         
  output [3:0]   ZQSFP_TXP,         
  output [3:0]   ZQSFP_TXN, 
  inout          QSFP_I2C_SCL,
  inout          QSFP_I2C_SDA,
  input          QSFP_MODPRSN,
  input          QSFP_INTN,
  output         QSFP_INITMODE,
  output         QSFP_MODSELN,
  output         QSFP_RESETN,
 
  //QSFPDD
  input  [7:0]   QSFPDD_RXP,         
  input  [7:0]   QSFPDD_RXN,         
  output [7:0]   QSFPDD_TXP,         
  output [7:0]   QSFPDD_TXN,  
  inout          QSFPDD_I2C_SCL,
  inout          QSFPDD_I2C_SDA,
  input          QSFPDD_MODPRSN,
  input          QSFPDD_INTN,
  output         QSFPDD_INITMODE,
  output         QSFPDD_MODSELN,
  output         QSFPDD_RESETN,   
  
 //PCIE
  input          PCIE_RC_PERSTN,
  input  [15:0]  PCIE_RC_RXP,         
  input  [15:0]  PCIE_RC_RXN,         
  output [15:0]  PCIE_RC_TXP,         
  output [15:0]  PCIE_RC_TXN, 
 
 //Ethernet
  output         ETH_RSTN,
  input          ETH_INTN, 
  inout          ETH_MDIO,
  output         ETH_MDC,  
  input          ETH_SGMII_RXN,
  input          ETH_SGMII_RXP,
  output         ETH_SGMII_TXN,
  output         ETH_SGMII_TXP,
  
 //Clock cleaner
  inout          CLKCLEANER_SCL,
  inout          CLKCLEANER_SDA,
  inout  [6:0]   CLKCLEANER_GPIO, 
  input  [1:0]   CLKCLEANER_STATUS, 
  output [1:0]   CLKCLEANER_INSEL0, 
  output [1:0]   CLKCLEANER_INSEL1, 
  output [1:0]   CLEARNER_RECOVERY_N, 
  output [1:0]   CLEARNER_RECOVERY_P,  
  input          CLEARNER_SYSTEM_N,
  input          CLEARNER_SYSTEM_P,
  
 //USB
  inout          USB_SCL,
  inout          USB_SDA,
  input          USB_RESETN,   
  input          USB_FPGA_CLK,
  output [1:0]   USB_ADDR, 
  inout  [7:0]   USB_DATA,  
  input          USB_WRN,
  input          USB_RDN,
  input          USB_OEN,
  output         USB_FULL,
  output         USB_EMPTY, 
 
 //Sodim 
  input          SODIMM_RZQ,
  input          SODIMM_REFCLKP,
  output         MEM_CLKN,
  output         MEM_CLKP,
  inout  [33:0]  MEM_DQA,   
  inout  [33:0]  MEM_DQB,   
  inout  [3:0]   MEM_DQSAN,
  inout  [3:0]   MEM_DQSAP,
  inout  [3:0]   MEM_DQSBN,
  inout  [3:0]   MEM_DQSBP,
  inout  [3:0]   MEM_DMAN,
  inout  [3:0]   MEM_DMBN,
  inout          MEM_DQS_ADDR_CMDN,
  inout          MEM_DQS_ADDR_CMDP,
  inout  [8:0]   MEM_DQ_ADDR_CMD,
  output [26:0]  MEM_ADDR_CMD,   
  input          MEM_ADDR_CMD27,
  output         MEM_ADDR_CMD28,
  output         MEM_ADDR_CMD29,
  output         MEM_ADDR_CMD30,
  
 //HPS   
  output         DDR4_COMP_CLKP,
  output         DDR4_COMP_CLKN,
  output [16:0]  DDR4_COMP_A,
  output         DDR4_COMP_ACTN,
  output [1:0]   DDR4_COMP_BA,
  output [1:0]   DDR4_COMP_BG,
  output         DDR4_COMP_CKE,
  output         DDR4_COMP_CSN,
  output         DDR4_COMP_ODT,
  output         DDR4_COMP_RESETN,
  output         DDR4_COMP_PAR,
  input          DDR4_COMP_ALERTN,
  input          DDR4_COMP_RZQ,
  input          DDR4_COMP_REFCLKP,
  inout [8:0]    DDR4_COMP_DBIN,
  inout [71:0]   DDR4_COMP_DQ,
  inout [8:0]    DDR4_COMP_DQSP,
  inout [8:0]    DDR4_COMP_DQSN,
  inout [47:0]   HPS_GPIO  
);

endmodule	