// ram1.v

// Generated using ACDS version 22.4 94

`timescale 1 ps / 1 ps
module ram1 (
		input  wire [31:0] data,    //    data.datain
		output wire [31:0] q,       //       q.dataout
		input  wire [9:0]  address, // address.address
		input  wire        wren,    //    wren.wren
		input  wire        clock,   //   clock.clk
		input  wire        aclr,    //    aclr.reset
		input  wire        rden     //    rden.rden
	);

	ram1_ram_1port_2010_evrarkq ram_1port_0 (
		.data    (data),    //   input,  width = 32,    data.datain
		.q       (q),       //  output,  width = 32,       q.dataout
		.address (address), //   input,  width = 10, address.address
		.wren    (wren),    //   input,   width = 1,    wren.wren
		.clock   (clock),   //   input,   width = 1,   clock.clk
		.aclr    (aclr),    //   input,   width = 1,    aclr.reset
		.rden    (rden)     //   input,   width = 1,    rden.rden
	);

endmodule
